`timescale 1ns/1ns
module JOYBUS_rx (
    input clk, rst_n,
    output [7:0] jb_cntlr_status,
    output [15:0] jb_cntlr_data,
);
    
endmodule